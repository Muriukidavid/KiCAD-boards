* opamp simulation
.include components.cir
XU1  3 6 5 4 2 OPAMP
R1  6 1 1K
R2  3 6 10K
V1  5 1 AC1
V2  3 5 AC2
XP1  2 5 4 PWR

.op
.tran 0.3m 1m 
.end
