* BJT characteristics

RB 1 2 1Meg
RC 4 3 1k	
Q1 3 2 0 BC107B 
V1 1 0 dc 12
V2 4 0 dc 10

.model BC107B   NPN(Is=7.049f Xti=3 Eg=1.11 Vaf=59.59 Bf=381.7 Ise=59.74f
+               Ne=1.522 Ikf=3.289 Nk=.5 Xtb=1.5 Br=2.359 Isc=192.9p Nc=1.954
+               Ikr=7.807 Rc=1.427 Cjc=5.38p Mjc=.329 Vjc=.6218 Fc=.5 Cje=11.5p
+               Mje=.2718 Vje=.5 Tr=10n Tf=438p Itf=5.716 Xtf=14.51 Vtf=10)
*       PHILIPS     pid=bc107b  case=TO18
*       91-08-02 dsq

.dc V2 0 10 0.1 V1 1.5 3.5 0.5 

************
.control
run
plot v(4,3)/1k vs v(3) 
.endc
************

.end
