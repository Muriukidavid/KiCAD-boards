* /home/karibe/src/kicad_boards/voltage_divider/voltage_divider.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 06 Jun 2017 10:51:29 AM EAT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R2  vout 0 10k		
R1  vout vin 3.9k		
v1  vin 0 DC 3.3		

.op
.tran 0.5s 1s
.tf v(vout,0) v1
.control
run
print all
*print dc v1#branch
*print vin
*print R2
.endc

*.control
*dc v1 3.3 3.3 0.1
*display
*.endc

.end
quit
