.title KiCad schematic
v1 0 vin DC 0 AC 1
R1 vout vin 1K
C1 vout 0 1.59uF
.ac dec 10 1 1Meg 
.control
run 
*Magnitude dB plot for vout on log scale 
plot vdb(vout) xlog 
*Phase degrees plot for vout on log scale 
plot {57.29*vp(vout)} xlog 
.endc
.end
