* /home/karibe/src/kicad_boards/BJT_amplifier/BJT_amplifier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 07 Jun 2017 01:32:35 AM EAT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  1 0 DC 12		
R1  2 1 1Meg		
R2  4 3 1k		
v2  4 0 DC 10		
Q1  3 2 0 BC107B		

.MODEL BJT1 NPN(BF=200 CJC=20pf CJE=20pf IS=1E16)

.model BC107B   NPN(Is=7.049f Xti=3 Eg=1.11 Vaf=59.59 Bf=381.7 Ise=59.74f
+               Ne=1.522 Ikf=3.289 Nk=.5 Xtb=1.5 Br=2.359 Isc=192.9p Nc=1.954
+               Ikr=7.807 Rc=1.427 Cjc=5.38p Mjc=.329 Vjc=.6218 Fc=.5 Cje=11.5p
+               Mje=.2718 Vje=.5 Tr=10n Tf=438p Itf=5.716 Xtf=14.51 Vtf=10)

.dc V2 0 10 0.1 V1 1.5 3.5 0.5 

************
.control
run
plot v(4,3)/1k vs v(3) 
.endc
************

.end

.end
