* Components and subcircuits for use in spicedemo.cir

.INCLUDE LMV981.MOD

*P1 2 5 4 PWR
*              + g -     
.subckt PWR 1 2 3
  Vneg 1 2 3.3V
  Vpos 2 3 3.3V
.ends PWR_IN

* XU1 3 6 5 4 2 OPAMP
*             o - + p n
.subckt OPAMP 1 2 3 8 4
  * PINOUT ORDER  1   3   6  2  4   5
  * PINOUT ORDER +IN -IN +V -V OUT NSD
  Xopamp 3 2 4 5 1 NSD LMV981
.ends OPAMP

* V1  5 1 AC1
*              s g
.subckt AC1 1 2
  Vmic 2 1 ac SIN(0 0.2 440)
ends AC1

* AC_2 3 5 vout
.subckt AC2 1 2
  Rwire 1 2 10ohm
ends AC2


